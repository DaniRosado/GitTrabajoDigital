package Estados_pkg is
    type estados is (SJug, ExtPied, IntrApuesta, ResRonda, FinJug);
end package;